package shared_pkg;
parameter DATA_W = 128;
parameter KEY_L = 128;
event valid_is_high;
endpackage